`ifndef __ROM_VH
`define __ROM_VH

`define ROM_SIZE 1024       // Todo: determine the rom size

`endif