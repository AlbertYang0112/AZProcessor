`ifndef __SPM_VH
`define __SPM_VH

`endif