`ifndef __SPM_VH
`define __SPM_VH

`define SPM_SIZE        16384
`define SPM_DEPTH       4096
`define SPM_ADDR_W      12
`define SPM_ADDR_BUS    11:0
`define SPM_ADDR_LOC    11:0

`endif