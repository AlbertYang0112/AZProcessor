`ifndef __ROM_VH
`define __ROM_VH

`define ROM_SIZE 8192
`define ROM_DEPTH 2048
`define ROM_ADDR_W 11
`define ROM_ADDR_BUS 10:0
`define ROM_ADDR_LOC 10:0

`endif