`ifndef __CPU_VH
`define __CPU_VH

`endif