`ifndef __CLOCK_VH
`define __CLOCK_VH

`define OSC_FREQ    50000000    // Todo: fill in the correct freq
`define CLOCK_DIV   0
`define CLOCK_FREQ  25000000

`endif