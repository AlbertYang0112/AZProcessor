`ifnedf __BUS_VH
`define __BUS_VH

`endif