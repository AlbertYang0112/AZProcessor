`ifndef __GPIO_VH
`define __GPIO_VH

`endif