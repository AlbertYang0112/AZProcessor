`ifndef __ISA_VH
`define __ISA_VH

`endif