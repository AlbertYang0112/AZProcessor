`include "nettype.vh"
`include "bus.vh"
`include "stddef.vh"

module bus(
    input wire                      clk,
    input wire                      reset_,
    input wire                      m0Req_,
    input wire                      m1Req_,
    input wire                      m2Req_,
    input wire                      m3Req_,
    output wire                     m0Grnt_,
    output wire                     m1Grnt_,
    output wire                     m2Grnt_,
    output wire                     m3Grnt_,
    input wire [`WORD_ADDR_BUS]     m0Addr,
    input wire [`WORD_ADDR_BUS]     m1Addr,
    input wire [`WORD_ADDR_BUS]     m2Addr,
    input wire [`WORD_ADDR_BUS]     m3Addr,
    input wire                      m0As_,
    input wire                      m1As_,
    input wire                      m2As_,
    input wire                      m3As_,
    input wire                      m0RW,
    input wire                      m1RW,
    input wire                      m2RW,
    input wire                      m3RW,
    input wire [`WORD_DATA_BUS]     m0Data,
    input wire [`WORD_DATA_BUS]     m1Data,
    input wire [`WORD_DATA_BUS]     m2Data,
    input wire [`WORD_DATA_BUS]     m3Data,
    output wire [`WORD_ADDR_BUS]    sAddr,
    output wire                     sAs_,
    output wire                     sRW,
    output wire [`WORD_DATA_BUS]    sData,
    output wire                     s0CS_,
    output wire                     s1CS_,
    output wire                     s2CS_,
    output wire                     s3CS_,
    output wire                     s4CS_,
    output wire                     s5CS_,
    output wire                     s6CS_,
    output wire                     s7CS_,
    (* KEEP = "{TRUE|FALSE |SOFT}" *)input wire [`WORD_DATA_BUS]     s0RdData,
    input wire [`WORD_DATA_BUS]     s1RdData,
    input wire [`WORD_DATA_BUS]     s2RdData,
    input wire [`WORD_DATA_BUS]     s3RdData,
    (* KEEP = "{TRUE|FALSE |SOFT}" *)input wire [`WORD_DATA_BUS]     s4RdData,
    input wire [`WORD_DATA_BUS]     s5RdData,
    input wire [`WORD_DATA_BUS]     s6RdData,
    input wire [`WORD_DATA_BUS]     s7RdData,
    input wire                      s0Rdy_,
    input wire                      s1Rdy_,
    input wire                      s2Rdy_,
    input wire                      s3Rdy_,
    input wire                      s4Rdy_,
    input wire                      s5Rdy_,
    input wire                      s6Rdy_,
    input wire                      s7Rdy_,
    output wire [`WORD_DATA_BUS]    mRdData,
    output wire                     mRdy_
);

    bus_arbiter BusArbiter(
        .clk(clk),
        .reset_(reset_),
        .m0Req_(m0Req_),
        .m1Req_(m1Req_),
        .m2Req_(m2Req_),
        .m3Req_(m3Req_),
        .m0Grnt_(m0Grnt_),
        .m1Grnt_(m1Grnt_),
        .m2Grnt_(m2Grnt_),
        .m3Grnt_(m3Grnt_)
    );
    
    bus_master_mux BusMasterMux(
        .m0Addr(m0Addr),
        .m1Addr(m1Addr),
        .m2Addr(m2Addr),
        .m3Addr(m3Addr),
        .m0As_(m0As_),
        .m1As_(m1As_),
        .m2As_(m2As_),
        .m3As_(m3As_),
        .m0RW(m0RW),
        .m1RW(m1RW),
        .m2RW(m2RW),
        .m3RW(m3RW),
        .m0Data(m0Data),
        .m1Data(m1Data),
        .m2Data(m2Data),
        .m3Data(m3Data),
        .m0Grnt_(m0Grnt_),
        .m1Grnt_(m1Grnt_),
        .m2Grnt_(m2Grnt_),
        .m3Grnt_(m3Grnt_),
        .sAddr(sAddr),
        .sAs_(sAs_),
        .sRW(sRW),
        .sData(sData)
    );

    bus_addr_dec BusAddrDec(
        .sAddr(sAddr),
        .s0CS_(s0CS_),
        .s1CS_(s1CS_),
        .s2CS_(s2CS_),
        .s3CS_(s3CS_),
        .s4CS_(s4CS_),
        .s5CS_(s5CS_),
        .s6CS_(s6CS_),
        .s7CS_(s7CS_)
    );

    bus_slave_mux BusSlaveMux(
        .s0CS_(s0CS_),
        .s1CS_(s1CS_),
        .s2CS_(s2CS_),
        .s3CS_(s3CS_),
        .s4CS_(s4CS_),
        .s5CS_(s5CS_),
        .s6CS_(s6CS_),
        .s7CS_(s7CS_),
        .s0RdData(s0RdData),
        .s1RdData(s1RdData),
        .s2RdData(s2RdData),
        .s3RdData(s3RdData),
        .s4RdData(s4RdData),
        .s5RdData(s5RdData),
        .s6RdData(s6RdData),
        .s7RdData(s7RdData),
        .s0Rdy_(s0Rdy_),
        .s1Rdy_(s1Rdy_),
        .s2Rdy_(s2Rdy_),
        .s3Rdy_(s3Rdy_),
        .s4Rdy_(s4Rdy_),
        .s5Rdy_(s5Rdy_),
        .s6Rdy_(s6Rdy_),
        .s7Rdy_(s7Rdy_),
        .mRdData(mRdData),
        .mRdy_(mRdy_)
    );


endmodule
