`ifnedf __ROM_VH
`define __ROM_VH

`endif