`ifndef __NETTYPE_H
`define __NETTYPE_H

`default_nettype none

`endif
