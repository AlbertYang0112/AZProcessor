
`define ENABLE 1
`define DISABLE 0
`define ASSERT 1
`define CLEAR 0