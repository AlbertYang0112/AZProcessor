`ifndef __GOLBAL_CONFIG_VH
`define __GOLBAL_CONFIG_VH

//`define POSITIVE_RESET NaN
`define NEGATIVE_RESET NaN
`define POSITIVE_MEMORY NaN
//`define NEGATIVE_MOMORY NaN
`define IMPLEMENT_TIMER NaN
`define IMPLEMENT_UART NaN
`define IMPLEMENT_GPIO NaN
`define RESET_EDGE negedge
`define RESET_ENABLE 1'b0
`define RESET_DISABLE 1'b1
`define MEM_ENABLE 1'b1
`define MEM_DISABLE 1'b0
`endif